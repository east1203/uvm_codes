`ifndef TEST__SV
`define TEST__SV

//program automatic test;
program test;

initial begin

  run_test("base_case");

end

endprogram

`endif
