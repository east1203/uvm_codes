
//`define RESULT_MON_PRINT
`define CMD_MON_PRINT
//`define MODEL_PRINT
