
package tb_pkg;
  import uvm_pkg::*;

  `include "uvm_macros.svh"

  `include "transaction.sv"
  `include "sequencer.sv"
  `include "driver.sv"
  `include "env.sv"
  `include "base_test.sv"
  `include "cases.sv"


endpackage


