

`ifndef PKG__SV
`define PKG__SV

package pkg;

`include "uvm_macros.svh"

import uvm_pkg::*;

`include  "transaction.sv"

endpackage


`endif





